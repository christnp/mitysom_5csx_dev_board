
module gbl_clock (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
